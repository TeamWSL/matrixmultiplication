`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 07/10/2024 09:03:53 AM
// Design Name: 
// Module Name: systolicarraytb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module tb_systolic_array_8x8;
    reg clk;
    reg reset;
    reg signed [7:0] A [0:3][0:3];
    reg signed [7:0] B [0:3][0:3];
    wire signed [15:0] C [0:3][0:3];

    matmul4x4 uut (
        .a(A),
        .b(B),
        .c(C)
    );

    initial begin

        // Initialize matrix A
        A[0][0] = 8'd1; A[0][1] = 8'd0; A[0][2] = 8'd0; A[0][3] = 8'd0; A[0][4] = 8'd0; A[0][5] = 8'd0; A[0][6] = 8'd0; A[0][7] = 8'd0;
        A[1][0] = 8'd0; A[1][1] = 8'd1; A[1][2] = 8'd0; A[1][3] = 8'd0; A[1][4] = 8'd0; A[1][5] = 8'd0; A[1][6] = 8'd0; A[1][7] = 8'd0;
        A[2][0] = 8'd0; A[2][1] = 8'd0; A[2][2] = 8'd1; A[2][3] = 8'd0; A[2][4] = 8'd0; A[2][5] = 8'd0; A[2][6] = 8'd0; A[2][7] = 8'd0;
        A[3][0] = 8'd0; A[3][1] = 8'd0; A[3][2] = 8'd0; A[3][3] = 8'd1; A[3][4] = 8'd0; A[3][5] = 8'd0; A[3][6] = 8'd0; A[3][7] = 8'd0;
        A[4][0] = 8'd0; A[4][1] = 8'd0; A[4][2] = 8'd0; A[4][3] = 8'd0; A[4][4] = 8'd1; A[4][5] = 8'd0; A[4][6] = 8'd0; A[4][7] = 8'd0;
        A[5][0] = 8'd0; A[5][1] = 8'd0; A[5][2] = 8'd0; A[5][3] = 8'd0; A[5][4] = 8'd0; A[5][5] = 8'd1; A[5][6] = 8'd0; A[5][7] = 8'd0;
        A[6][0] = 8'd0; A[6][1] = 8'd0; A[6][2] = 8'd0; A[6][3] = 8'd0; A[6][4] = 8'd0; A[6][5] = 8'd0; A[6][6] = 8'd1; A[6][7] = 8'd0;
        A[7][0] = 8'd0; A[7][1] = 8'd0; A[7][2] = 8'd0; A[7][3] = 8'd0; A[7][4] = 8'd0; A[7][5] = 8'd0; A[7][6] = 8'd0; A[7][7] = 8'd1;
        

        // Initialize matrix B
        B[0][0] = 8'd1; B[0][1] = 8'd2; B[0][2] = 8'd3; B[0][3] = 8'd4; B[0][4] = 8'd5; B[0][5] = 8'd6; B[0][6] = 8'd7; B[0][7] = 8'd8;
        B[1][0] = 8'd9; B[1][1] = 8'd10; B[1][2] = 8'd11; B[1][3] = 8'd12; B[1][4] = 8'd13; B[1][5] = 8'd14; B[1][6] = 8'd15; B[1][7] = 8'd16;
        B[2][0] = 8'd17; B[2][1] = 8'd18; B[2][2] = 8'd19; B[2][3] = 8'd20; B[2][4] = 8'd21; B[2][5] = 8'd22; B[2][6] = 8'd23; B[2][7] = 8'd24;
        B[3][0] = 8'd25; B[3][1] = 8'd26; B[3][2] = 8'd27; B[3][3] = 8'd28; B[3][4] = 8'd29; B[3][5] = 8'd30; B[3][6] = 8'd31; B[3][7] = 8'd32;
        B[4][0] = 8'd33; B[4][1] = 8'd34; B[4][2] = 8'd35; B[4][3] = 8'd36; B[4][4] = 8'd37; B[4][5] = 8'd38; B[4][6] = 8'd39; B[4][7] = 8'd40;
        B[5][0] = 8'd41; B[5][1] = 8'd42; B[5][2] = 8'd43; B[5][3] = 8'd44; B[5][4] = 8'd45; B[5][5] = 8'd46; B[5][6] = 8'd47; B[5][7] = 8'd48;
        B[6][0] = 8'd49; B[6][1] = 8'd50; B[6][2] = 8'd51; B[6][3] = 8'd52; B[6][4] = 8'd53; B[6][5] = 8'd54; B[6][6] = 8'd55; B[6][7] = 8'd56;
        B[7][0] = 8'd57; B[7][1] = 8'd58; B[7][2] = 8'd59; B[7][3] = 8'd60; B[7][4] = 8'd61; B[7][5] = 8'd62; B[7][6] = 8'd63; B[7][7] = 8'd64;

        #100;

        // Display the result matrix C
        $display("Matrix C:");
        for (integer i = 0; i < 8; i = i + 1) begin
            $display("%d %d %d %d %d %d %d %d",
                C[i][0], C[i][1], C[i][2], C[i][3],
                C[i][4], C[i][5], C[i][6], C[i][7]);
        end

    end

endmodule



