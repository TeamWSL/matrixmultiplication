`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 07/11/2024 07:31:28 PM
// Design Name: 
// Module Name: matmul4x4
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module matmul4x4(
    input wire signed [7:0] a [0:3][0:3],
    input wire signed [7:0] b [0:3][0:3],
    output reg signed [15:0] c [0:3][0:3]
    );
    pematmul pm1(.a1(a[0][3]), .b1(b[3][0]), .a2(a[0][2]), .b2(b[2][0]), .a3(a[0][1]), .b3(b[1][0]), .a4(a[0][0]), .b4(b[0][0]), .c(c[0][0]));
    pematmul pm2(.a1(a[0][3]), .b1(b[3][1]), .a2(a[0][2]), .b2(b[2][1]), .a3(a[0][1]), .b3(b[1][1]), .a4(a[0][0]), .b4(b[0][1]), .c(c[0][1]));
    pematmul pm3(.a1(a[0][3]), .b1(b[3][2]), .a2(a[0][2]), .b2(b[2][2]), .a3(a[0][1]), .b3(b[1][2]), .a4(a[0][0]), .b4(b[0][2]), .c(c[0][2]));
    pematmul pm4(.a1(a[0][3]), .b1(b[3][3]), .a2(a[0][2]), .b2(b[2][3]), .a3(a[0][1]), .b3(b[1][3]), .a4(a[0][0]), .b4(b[0][3]), .c(c[0][3]));
    pematmul pm5(.a1(a[1][3]), .b1(b[3][0]), .a2(a[1][2]), .b2(b[2][0]), .a3(a[1][1]), .b3(b[1][0]), .a4(a[1][0]), .b4(b[0][0]), .c(c[1][0]));
    pematmul pm6(.a1(a[1][3]), .b1(b[3][1]), .a2(a[1][2]), .b2(b[2][1]), .a3(a[1][1]), .b3(b[1][1]), .a4(a[1][0]), .b4(b[0][1]), .c(c[1][1]));
    pematmul pm7(.a1(a[1][3]), .b1(b[3][2]), .a2(a[1][2]), .b2(b[2][2]), .a3(a[1][1]), .b3(b[1][2]), .a4(a[1][0]), .b4(b[0][2]), .c(c[1][2]));
    pematmul pm8(.a1(a[1][3]), .b1(b[3][3]), .a2(a[1][2]), .b2(b[2][3]), .a3(a[1][1]), .b3(b[1][3]), .a4(a[1][0]), .b4(b[0][3]), .c(c[1][3]));
    pematmul pm9(.a1(a[2][3]), .b1(b[3][0]), .a2(a[2][2]), .b2(b[2][0]), .a3(a[2][1]), .b3(b[1][0]), .a4(a[2][0]), .b4(b[0][0]), .c(c[2][0]));
    pematmul pm10(.a1(a[2][3]), .b1(b[3][1]), .a2(a[2][2]), .b2(b[2][1]), .a3(a[2][1]), .b3(b[1][1]), .a4(a[2][0]), .b4(b[0][1]), .c(c[2][1]));
    pematmul pm11(.a1(a[2][3]), .b1(b[3][2]), .a2(a[2][2]), .b2(b[2][2]), .a3(a[2][1]), .b3(b[1][2]), .a4(a[2][0]), .b4(b[0][2]), .c(c[2][2]));
    pematmul pm12(.a1(a[2][3]), .b1(b[3][3]), .a2(a[2][2]), .b2(b[2][3]), .a3(a[2][1]), .b3(b[1][3]), .a4(a[2][0]), .b4(b[0][3]), .c(c[2][3]));
    pematmul pm13(.a1(a[3][3]), .b1(b[3][0]), .a2(a[3][2]), .b2(b[2][0]), .a3(a[3][1]), .b3(b[1][0]), .a4(a[3][0]), .b4(b[0][0]), .c(c[3][0]));
    pematmul pm14(.a1(a[3][3]), .b1(b[3][1]), .a2(a[3][2]), .b2(b[2][1]), .a3(a[3][1]), .b3(b[1][1]), .a4(a[3][0]), .b4(b[0][1]), .c(c[3][1]));
    pematmul pm15(.a1(a[3][3]), .b1(b[3][2]), .a2(a[3][2]), .b2(b[2][2]), .a3(a[3][1]), .b3(b[1][2]), .a4(a[3][0]), .b4(b[0][2]), .c(c[3][2]));
    pematmul pm16(.a1(a[3][3]), .b1(b[3][3]), .a2(a[3][2]), .b2(b[2][3]), .a3(a[3][1]), .b3(b[1][3]), .a4(a[3][0]), .b4(b[0][3]), .c(c[3][3]));
endmodule
